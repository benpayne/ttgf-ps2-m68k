`default_nettype none
`timescale 1ns / 1ps

/* This testbench just instantiates the module and makes some convenient wires
   that can be driven / tested by the cocotb test.py.
*/
module tb ();

  // Dump the signals to a VCD file. You can view it with gtkwave.
  initial begin
    $dumpfile("tb.vcd");
    $dumpvars(0, tb);
    #1;
  end

  // Wire up the inputs and outputs:
  reg clk;
  reg rst_n;
  reg ena;
  reg [7:0] ui_in;
  reg [7:0] uio_in;
  wire [7:0] uo_out;
  wire [7:0] uio_out;
  wire [7:0] uio_oe;

  // Power supply wires for GF180
  wire VPWR;
  wire VGND;
  assign VPWR = 1'b1;
  assign VGND = 1'b0;

  wire ps2_clk;
  wire ps2_data;
  wire clear_int;
  wire valid;
  wire interupt;
  wire cs;
  wire data_rdy;
  wire fifo_full;

  assign ui_in[0] = ps2_clk;
  assign ui_in[1] = ps2_data;
  assign ui_in[2] = clear_int;
  assign ui_in[3] = cs;

  assign valid = uo_out[0];
  assign interupt = uo_out[1];
  assign data_rdy = uo_out[2];
  assign fifo_full = uo_out[3];

  // Replace tt_um_example with your module name:
  tt_um_benpayne_ps2_decoder user_project (

      // Include power ports (required for GF180):
      .VPWR(VPWR),
      .VGND(VGND),

      .clk    (clk),      // clock
      .ena    (ena),      // enable - goes high when design is selected
      .rst_n  (rst_n),    // not reset
      .ui_in  (ui_in),    // Dedicated inputs
      .uio_in (uio_in),   // IOs: Input path
      .uio_oe (uio_oe),   // IOs: Enable path (active high: 0=input, 1=output)
      .uio_out(uio_out),  // IOs: Output path
      .uo_out (uo_out)    // Dedicated outputs
  );

endmodule
